library verilog;
use verilog.vl_types.all;
entity ProcessorMIPS_vlg_vec_tst is
end ProcessorMIPS_vlg_vec_tst;
